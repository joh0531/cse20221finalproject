module obstacle_DE2 (
	input CLOCK_50, // 50 MHz
	input [0:0] KEY,
	output VGA_CLK, // VGA Clock
	output VGA_HS, // VGA H_SYNC
	output VGA_VS, // VGA V_SYNC
	output VGA_BLANK, // VGA BLANK
	output VGA_SYNC, // VGA SYNC
	output [9:0] VGA_R, // VGA Red[9:0]
	output [9:0] VGA_G, // VGA Green[9:0]
	output [9:0] VGA_B // VGA Blue[9:0]
	);
	
	wire [2:0] color;
	wire [7:0] x;
	wire [6:0] y;
	wire plot;
	
	processor (
	.clk (CLOCK_50),
	.reset (~KEY[0]),
	.xpos (x),
	.ypos (y),
	.color (color),
	.plot (plot)
	);
	
	vga_adapter VGA(
	.resetn(KEY[0]),
	.clock(CLOCK_50),
	.colour(color),
	.x(x),
	.y(y),
	.plot(plot),
	/* Signals for the DAC to drive the monitor. */
	.VGA_R(VGA_R),
	.VGA_G(VGA_G),
	.VGA_B(VGA_B),
	.VGA_HS(VGA_HS),
	.VGA_VS(VGA_VS),
	.VGA_BLANK(VGA_BLANK),
	.VGA_SYNC(VGA_SYNC),
	.VGA_CLK(VGA_CLK)
	);
	
	defparam VGA.RESOLUTION = "160x120";
	defparam VGA.MONOCHROME = "FALSE";
	defparam VGA.BITS_PER_COLOUR_CHANNEL = 1;
	defparam VGA.BACKGROUND_IMAGE = "obstacle_course.mif";
	
endmodule